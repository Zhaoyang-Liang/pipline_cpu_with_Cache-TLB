`timescale 1ns / 1ps
//*************************************************************************
//   > �ļ���: wb.v
//   > ����  :�弶��ˮCPU��д��ģ��
//   > ����  : LOONGSON
//   > ����  : 2016-04-14
//*************************************************************************
module wb(                       // д�ؼ�
    input          WB_valid,     // д�ؼ���Ч
    input  [155:0] MEM_WB_bus_r, // MEM->WB����
    output         rf_wen,       // �Ĵ���дʹ��
    output [  4:0] rf_wdest,     // �Ĵ���д��ַ
    output [ 31:0] rf_wdata,     // �Ĵ���д����
    output         WB_over,      // WBģ��ִ�����

     //5����ˮ�����ӿ�
    input             clk,       // ʱ��
    input             resetn,    // ��λ�źţ��͵�ƽ��Ч
    output [ 32:0] exc_bus,      // Exception pc����
    output [  4:0] WB_wdest,     // WB��Ҫд�ؼĴ����ѵ�Ŀ���ַ��
    output         cancel,       // syscall��eret����д�ؼ�ʱ�ᷢ��cancel�źţ�
                                  // ȡ���Ѿ�ȡ��������������ˮ��ִ�е�ָ��
 
    // ������·�������
    output     [ 31:0] WB_result,   // WB�������������·

     //չʾPC��HI/LOֵ
    output [ 31:0] WB_pc,
    output [ 31:0] HI_data,
    output [ 31:0] LO_data,

    // �۲�CP0�Ĵ��������ڵ���/��ʾ��
    output [ 31:0] cp0_status,
    output [ 31:0] cp0_cause,
    output [ 31:0] cp0_epc
);
//-----{MEM->WB����}begin    
    //MEM������result
    wire [31:0] mem_result;
    //HI/LO����
    wire [31:0] lo_result;
    wire        hi_write;
    wire        lo_write;
    
    //�Ĵ�����дʹ�ܺ�д��ַ
    wire wen;
    wire [4:0] wdest;
    
    //д����Ҫ�õ�����Ϣ
    wire mfhi;
    wire mflo;
    wire mtc0;
    wire mfc0;
    wire [7 :0] cp0r_addr;
    wire       syscall;   //syscall��eret��д�ؼ�������Ĳ��� 
    wire       eret;
    
    //pc
    wire [31:0] pc;    
    wire        mem_ex_adel_wb;
    wire        mem_ex_ades_wb;
    wire        mem_ex_tlbl_wb;
    wire        mem_ex_tlbs_wb;
    wire        mem_ex_mod_wb;
    wire [31:0] mem_badvaddr_wb;
    wire        brk_wb;
    assign {wen,
            wdest,
            mem_result,
            lo_result,
            hi_write,
            lo_write,
            mfhi,
            mflo,
            mtc0,
            mfc0,
            cp0r_addr,
            syscall,
            brk_wb,
            eret,
            mem_ex_adel_wb,
            mem_ex_ades_wb,
            mem_ex_tlbl_wb,
            mem_ex_tlbs_wb,
            mem_ex_mod_wb,
            mem_badvaddr_wb,
            pc} = MEM_WB_bus_r;
//-----{MEM->WB����}end

//-----{HI/LO�Ĵ���}begin
    //HI���ڴ�ų˷�����ĸ�32λ
    //LO���ڴ�ų˷�����ĵ�32λ
    reg [31:0] hi;
    reg [31:0] lo;
    
    //Ҫд��HI�����ݴ����mem_result��
    always @(posedge clk)
    begin
        if (hi_write)
        begin
            hi <= mem_result;
        end
    end
    //Ҫд��LO�����ݴ����lo_result��
    always @(posedge clk)
    begin
        if (lo_write)
        begin
            lo <= lo_result;
        end
    end
//-----{HI/LO�Ĵ���}end


// //-----{cp0�Ĵ���}begin
// // cp0�Ĵ�������Э������0�Ĵ���
// // ����Ŀǰ��Ƶ�CPU�����걸�����õ���cp0�Ĵ���Ҳ����
// // ����ʱֻʵ��STATUS(12.0),CAUSE(13.0),EPC(14.0)������
// // ÿ��CP0�Ĵ�������ʹ��5λ��cp0��
//    wire [31:0] cp0r_status;
//    wire [31:0] cp0r_cause;
//    wire [31:0] cp0r_epc;
   
//    //дʹ��
//    wire status_wen;
//    //wire cause_wen;
//    wire epc_wen;
//    assign status_wen = mtc0 & (cp0r_addr=={5'd12,3'd0});
//    assign epc_wen    = mtc0 & (cp0r_addr=={5'd14,3'd0});
   
//    //cp0�Ĵ�����
//    wire [31:0] cp0r_rdata;
//    assign cp0r_rdata = (cp0r_addr=={5'd12,3'd0}) ? cp0r_status :
//                        (cp0r_addr=={5'd13,3'd0}) ? cp0r_cause  :
//                        (cp0r_addr=={5'd14,3'd0}) ? cp0r_epc : 32'd0;
   
//    //STATUS�Ĵ���
//    //Ŀǰֻʵ��STATUS[1]λ����EXL��
//    //EXL��Ϊ����ɶ�д������Ҫstatu_wen
//    reg status_exl_r;
//    assign cp0r_status = {30'd0,status_exl_r,1'b0};
//    always @(posedge clk)
//    begin
//        if (!resetn || eret)
//        begin
//            status_exl_r <= 1'b0;
//        end
//        else if (syscall)
//        begin
//            status_exl_r <= 1'b1;
//        end
//        else if (status_wen)
//        begin
//            status_exl_r <= mem_result[1];
//        end
//    end
   
//    //CAUSE�Ĵ���
//    //Ŀǰֻʵ��CAUSE[6:2]λ����ExcCode��,���Exception����
//    //ExcCode��Ϊ���ֻ��������д���ʲ���Ҫcause_wen
//    reg [4:0] cause_exc_code_r;
//    assign cp0r_cause = {25'd0,cause_exc_code_r,2'd0};
//    always @(posedge clk)
//    begin
//        if (syscall)
//        begin
//            cause_exc_code_r <= 5'd8;
//        end
//    end
   
//    //EPC�Ĵ���
//    //��Ų�������ĵ�ַ
//    //EPC������Ϊ����ɶ�д�ģ�����Ҫepc_wen
//    reg [31:0] epc_r;
//    assign cp0r_epc = epc_r;
//    always @(posedge clk)
//    begin
//        if (syscall)
//        begin
//            epc_r <= pc;
//        end
//        else if (epc_wen)
//        begin
//            epc_r <= mem_result;
//        end
//    end
   
//    //syscall��eret������cancel�ź�
//    assign cancel = (syscall | eret) & WB_over;
// //-----{cp0�Ĵ���}begin

//-----{CP0ģ��ʵ����}begin-----
   // CP0�Ĵ���������
   wire [31:0] cp0r_rdata;
   // CP0�Ĵ���ֵ�������쳣����
   wire [31:0] cp0r_status;
   wire [31:0] cp0r_cause;
   wire [31:0] cp0r_epc;
   // CP0������쳣�����ź�
   wire        cp0_cancel;
   wire        cp0_exc_valid;
   wire [31:0] cp0_exc_pc;
   wire        cp0_int;      // CP0�ж��ź�
   
   // ͳһ�쳣�����ź���������������ʹ�ã�
   wire        wb_ex_valid;
   wire [4:0]  wb_ex_code;
   wire        wb_ex_bd;
   wire [31:0] wb_ex_pc;
   wire        wb_badvaddr_valid;
   wire [31:0] wb_badvaddr;
   
   // �쳣�ٲ��߼������ȼ����ж� > ��ַ�� > BREAK > SYSCALL��
   // ע�⣺�ж���CP0ģ���⣬ͨ��c0_int�źŴ���
   // ����cp0_int��CP0ʵ������ſ��ã������ȼ�����ж��쳣��Ȼ����CP0ʵ������ϲ��ж�
   assign wb_badvaddr_valid   = (mem_ex_tlbl_wb | mem_ex_tlbs_wb | mem_ex_mod_wb |
                                  mem_ex_adel_wb | mem_ex_ades_wb);
   assign wb_badvaddr         = mem_badvaddr_wb;
   
   // ���ж��쳣����ַ��BREAK��SYSCALL��
   wire        wb_ex_valid_no_int;
   wire [4:0]  wb_ex_code_no_int;
   assign wb_ex_valid_no_int  = (mem_ex_tlbl_wb | mem_ex_tlbs_wb | mem_ex_mod_wb |
                                mem_ex_adel_wb | mem_ex_ades_wb | brk_wb | syscall) ? WB_valid : 1'b0;
   assign wb_ex_code_no_int    = mem_ex_tlbl_wb ? 5'd2 :
                                mem_ex_tlbs_wb ? 5'd3 :
                                mem_ex_mod_wb  ? 5'd1 :
                                mem_ex_adel_wb ? 5'd4 :
                                mem_ex_ades_wb ? 5'd5 :
                                brk_wb ? 5'd9 :
                                5'd8; // SYSCALL

   always @(posedge clk) begin
       if (wb_ex_valid) begin
           $display("WB_EXC_ARB: code=%0d badvaddr=%h pc=%h", wb_ex_code, wb_badvaddr, pc);
       end
   end
   
   cp0 cp0_module(
       .clk         (clk         ),  // I, 1
       .resetn      (resetn      ),  // I, 1
       .mtc0        (mtc0        ),  // I, 1
       .mfc0        (mfc0        ),  // I, 1
       .cp0r_addr   (cp0r_addr   ),  // I, 8
       .wdata       (mem_result  ),  // I, 32
       .syscall     (syscall     ),  // I, 1
       .eret        (eret        ),  // I, 1
       .pc          (pc          ),  // I, 32
       .wb_valid    (WB_valid    ),  // I, 1
       .wb_over     (WB_over     ),  // I, 1
       // ͳһ�쳣����
       .ex_valid_i        (wb_ex_valid       ), // I, 1
       .ex_code_i         (wb_ex_code        ), // I, 5
       .ex_bd_i           (wb_ex_bd          ), // I, 1
       .ex_pc_i           (wb_ex_pc          ), // I, 32
       .badvaddr_valid_i  (wb_badvaddr_valid ), // I, 1
       .badvaddr_i        (wb_badvaddr       ), // I, 32
       .cp0r_rdata  (cp0r_rdata  ),  // O, 32
       .cancel      (cp0_cancel  ),  // O, 1
       .exc_valid   (cp0_exc_valid), // O, 1
       .exc_pc      (cp0_exc_pc  ),  // O, 32
       .cp0r_status (cp0r_status ),  // O, 32
       .cp0r_cause  (cp0r_cause  ),  // O, 32
       .cp0r_epc    (cp0r_epc    ),  // O, 32
       .c0_int      (cp0_int     )   // O, 1  // �ж��ź�
   );
   
   // ��CP0��cancel�ź����ӵ�WB��cancel���
   assign cancel = cp0_cancel;
   
   // �����쳣�ٲã������жϣ��ж����ȼ���ߣ�
   // ע�⣺cp0_int�����ѿ��ã�CP0ģ����ʵ������
   // wb_ex_valid_no_int�Ѿ�������WB_valid����������ֻ��Ҫ����cp0_int�����
   assign wb_ex_valid = (cp0_int && WB_valid) | wb_ex_valid_no_int;
   assign wb_ex_code  = cp0_int ? 5'd0 : wb_ex_code_no_int;  // �ж��쳣��Ϊ0
   assign wb_ex_bd    = 1'b0;       // �ӳٲۺ�������
   assign wb_ex_pc    = pc;         // �쳣PC����ַ����syscall��ȡ��ǰpc��
//-----{CP0ģ��ʵ����}end-----

//-----{WBִ�����}begin
    //WBģ�����в���������һ�������
    //��WB_valid����WB_over�ź�
    assign WB_over = WB_valid;
//-----{WBִ�����}end

//-----{WB->regfile�ź�}begin
    assign rf_wen   = wen & WB_over;
    assign rf_wdest = wdest;
    assign rf_wdata = mfhi ? hi :
                      mflo ? lo :
                      mfc0 ? cp0r_rdata : mem_result;

    assign WB_result = rf_wdata;  // ! ��·���
//-----{WB->regfile�ź�}end


//-----{Exception pc�ź�}begin-----
    // �쳣���ߣ�{�쳣��Ч�ź�, �쳣PC��ַ}
    // �쳣�����߼��ѷ�װ��CP0ģ����
    assign exc_bus = {cp0_exc_valid, cp0_exc_pc};
//-----{Exception pc�ź�}end-----

//-----{WBģ���destֵ}begin
   //ֻ����WBģ����Чʱ����д��Ŀ�ļĴ����Ų�������
    assign WB_wdest = rf_wdest & {5{WB_valid}};
//-----{WBģ���destֵ}end

//-----{չʾWBģ���PCֵ��HI/LO�Ĵ�����ֵ}begin
    assign WB_pc = pc;
    assign HI_data = hi;
    assign LO_data = lo;
//-----{չʾWBģ���PCֵ��HI/LO�Ĵ�����ֵ}end

//-----{����CP0�Ĵ������ڹ۲�}begin
    assign cp0_status = cp0r_status;
    assign cp0_cause  = cp0r_cause;
    assign cp0_epc    = cp0r_epc;
//-----{����CP0�Ĵ������ڹ۲�}end
endmodule

