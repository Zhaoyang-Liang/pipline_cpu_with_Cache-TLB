`timescale 1ns / 1ps
//*************************************************************************
//   > �ļ���: cp0.v
//   > ����  :Э������0��CP0��ģ�飬����ϵͳ���ƺ��쳣����
//   > ����  : 
//   > ����  : 
//*************************************************************************

`define EXC_ENTER_ADDR 32'd0     // Exception��ڵ�ַ���˴�ʵ�ֵ�Exceptionֻ��SYSCALL

module cp0(
    input             clk,       // ʱ��
    input             resetn,    // ��λ�źţ��͵�ƽ��Ч
    
    // ����WB���Ŀ����ź�
    input             mtc0,      // MTC0ָ���ʶ
    input             mfc0,      // MFC0ָ���ʶ
    input      [ 7:0] cp0r_addr, // CP0�Ĵ�����ַ {�Ĵ�����[4:0], ѡ����[2:0]}
    input      [31:0] wdata,     // д��CP0�����ݣ�����mem_result��
    
    // �쳣����ź�
    input             syscall,   // SYSCALLָ���ʶ
    input             eret,      // ERETָ���ʶ
    input      [31:0] pc,        // ��ǰPCֵ�����ڱ��浽EPC��
    input             wb_valid,  // WB����Ч�ź�
    input             wb_over,   // WB������ź�

    // ͳһ�쳣���ߣ�����WB�����ղþ���
    input             ex_valid_i,        // �쳣��Ч
    input      [ 4:0] ex_code_i,         // �쳣����
    input             ex_bd_i,           // �ӳٲ��쳣
    input      [31:0] ex_pc_i,           // �����쳣��PC����bd=1��Ϊ��֧PC��
    input             badvaddr_valid_i,  // �����ַ��Ч
    input      [31:0] badvaddr_i,        // �����ַ
    
    // CP0�Ĵ������������
    output     [31:0] cp0r_rdata,// CP0�Ĵ��������ݣ�����MFC0��
    
    // �쳣�������
    output            cancel,    // ȡ����ˮ���ź�
    output            exc_valid, // �쳣��Ч�ź�
    output     [31:0] exc_pc,    // �쳣��ڵ�ַ��ERET���ص�ַ
    
    // �Ĵ���ֵ����������쳣����
    output     [31:0] cp0r_status,// STATUS�Ĵ���ֵ
    output     [31:0] cp0r_cause, // CAUSE�Ĵ���ֵ
    output     [31:0] cp0r_epc,   // EPC�Ĵ���ֵ
    
    // �ж����
    output            c0_int      // �ж���Ч�ź�
);

// ��ַ���루reg_num[4:0], sel[2:0]��
wire [4:0] cp0_reg_num = cp0r_addr[7:3];
wire [2:0] cp0_sel     = cp0r_addr[2:0];
wire sel_status = (cp0_reg_num==5'd12) && (cp0_sel==3'd0);
wire sel_cause  = (cp0_reg_num==5'd13) && (cp0_sel==3'd0);
wire sel_epc    = (cp0_reg_num==5'd14) && (cp0_sel==3'd0);
wire sel_count  = (cp0_reg_num==5'd9)  && (cp0_sel==3'd0);   // COUNT�Ĵ���
wire sel_compare= (cp0_reg_num==5'd11) && (cp0_sel==3'd0);   // COMPARE�Ĵ���
wire sel_badvaddr = (cp0_reg_num==5'd8) && (cp0_sel==3'd0);  // BADVADDR�Ĵ���

// CP0�Ĵ�����status/cause/epc/badvaddr/count/compare
reg [31:0] status;
reg [31:0] cause;
reg [31:0] epc;
reg [31:0] badvaddr;
reg [31:0] count;      // COUNT�Ĵ�������ʱ��������
reg [31:0] compare;    // COMPARE�Ĵ�������ʱ���Ƚ�ֵ��

// STATUS�Ĵ���λ��
wire status_ie;        // bit 0: ȫ���ж�ʹ��
wire status_exl;       // bit 1: �쳣����
wire [7:0] status_im;  // bit 15:8: �ж�����λ

// CAUSE�Ĵ���λ��
wire cause_bd;         // bit 31: �ӳٲ۱�־
wire cause_ti;         // bit 30: ��ʱ���жϱ�־
wire [7:0] cause_ip;   // bit 15:8: �жϹ���λ
wire [4:0] cause_excode; // bit 6:2: �쳣����

// ��ʱ������ź�
reg time_tick;         // ��ʱ��ʱ�ӷ�Ƶ��ÿ����ʱ�����ڷ�תһ�Σ�
wire count_eq_compare; // COUNT == COMPARE
reg cause_ti_reg;     // ��ʱ���жϱ�־�Ĵ���

// STATUS��CAUSE�Ĵ���λ��ֵ
assign status_ie  = status[0];
assign status_exl = status[1];
assign status_im  = status[15:8];

assign cause_bd     = cause[31];
assign cause_ti     = cause[30];
assign cause_ip     = cause[15:8];
assign cause_excode = cause[6:2];

// ���� output: cp0r_status, cp0r_cause, cp0r_epc
assign cp0r_status = status;
assign cp0r_cause  = cause;
assign cp0r_epc    = epc;

// COUNT == COMPARE���
assign count_eq_compare = (count == compare);

// д�����ź�
wire status_wen;
wire cause_wen;
wire epc_wen;
wire count_wen;
wire compare_wen;
wire badvaddr_wen;
wire mtc0_wr;  // MTC0дʹ�ܣ��ų��쳣ʱд�룩

assign mtc0_wr      = mtc0 && wb_valid && !ex_valid_i; // �쳣ʱ��д��
assign status_wen   = mtc0_wr && sel_status;
assign cause_wen    = mtc0_wr && sel_cause;
assign epc_wen      = mtc0_wr && sel_epc;
assign count_wen    = mtc0_wr && sel_count;
assign compare_wen  = mtc0_wr && sel_compare;
assign badvaddr_wen = mtc0_wr && sel_badvaddr;

// STATUS�Ĵ���д���루֧��IE��EXL��IMλ��
wire [31:0] STATUS_WMASK;
assign STATUS_WMASK = 32'h0000_8103; // bit 0(IE), bit 1(EXL), bit 15:8(IM)

// CAUSE�Ĵ���д���루֧��IP[1:0]λ��
wire [31:0] CAUSE_WMASK;
assign CAUSE_WMASK = 32'h0000_0300;  // bit 9:8(IP[1:0])

// ��ʱ��ʱ�ӷ�Ƶ��ÿ����ʱ�����ڷ�תһ�Σ����ͼ���Ƶ�ʣ�
always @(posedge clk) begin
    if (!resetn) begin
        time_tick <= 1'b0;
    end else begin
        time_tick <= ~time_tick;
    end
end

// COUNT�Ĵ�������д����ÿ����ʱ����������
always @(posedge clk) begin
    if (!resetn) begin
        count <= 32'd0;
    end else begin
        if (count_wen) begin
            count <= wdata;
        end else if (time_tick) begin
            count <= count + 1'b1;
        end
    end
end

// COMPARE�Ĵ�������д��д��ʱ�����ʱ���ж�
always @(posedge clk) begin
    if (!resetn) begin
        compare <= 32'd0;
    end else begin
        if (compare_wen) begin
            compare <= wdata;
        end
    end
end

// ��ʱ���жϱ�־��cause_ti_reg��
always @(posedge clk) begin
    if (!resetn) begin
        cause_ti_reg <= 1'b0;
    end else begin
        if (compare_wen) begin
            cause_ti_reg <= 1'b0;  // д��COMPAREʱ���
        end else if (count_eq_compare) begin
            cause_ti_reg <= 1'b1;   // COUNT == COMPAREʱ��λ
        end
    end
end

// CP0�Ĵ������߼�
always @(posedge clk) begin
    if (!resetn) begin
        status <= 32'd0;
        cause  <= 32'd0;
        epc    <= 32'd0;
        badvaddr <= 32'd0;
    end else begin
        // MTC0д��
        if (status_wen) begin
            status <= (status & ~STATUS_WMASK) | (wdata & STATUS_WMASK);
        end
        if (cause_wen) begin
            cause <= (cause & ~CAUSE_WMASK) | (wdata & CAUSE_WMASK);
        end
        if (epc_wen) begin
            epc <= wdata;
        end
        if (badvaddr_wen) begin
            badvaddr <= wdata;
        end

        // ͳһ�쳣���������쳣��ͨ��ex_valid_i����
        // ע�⣺��Ϊ�ӳٲ��쳣ʱ��EPC��д��ָ֧��PC���� ex_pc_i��������ʱ������������Ƿ�+4
        if (ex_valid_i && wb_valid) begin
            status[1] <= 1'b1;                     // EXL
            cause[31] <= ex_bd_i;                  // BD
            cause[6:2] <= ex_code_i;               // ExcCode
            epc <= ex_bd_i ? ex_pc_i : ex_pc_i;   // ����д���֧PC�����PC
            if (badvaddr_valid_i) begin
                badvaddr <= badvaddr_i;
            end
        end
        
        // ERETָ����EXLλ
        if (eret && wb_valid) begin
            status[1] <= 1'b0;   // ��EXL
        end
        
        // CAUSE�Ĵ���λ����£��������£������쳣����Ӱ�죩
        // cause[30]: TIλ����ʱ���жϱ�־��
        if (!ex_valid_i || !wb_valid) begin
            cause[30] <= cause_ti_reg;
        end
        
        // cause[15:8]: IPλ���жϹ���λ��
        // IP[7] = TI����ʱ���жϣ�
        // IP[6:2] = �ⲿ�жϣ���δʵ�֣�����Ϊ0��
        // IP[1:0] = �����д����MTC0���ƣ�
        if (!ex_valid_i || !wb_valid) begin
            cause[15:8] <= {cause_ti_reg, 5'd0, cause[9:8]};
        end
    end
end

// MFC0��
assign cp0r_rdata = sel_status  ? status   :
                    sel_cause   ? cause    :
                    sel_epc     ? epc      :
                    sel_count   ? count    :
                    sel_compare ? compare  :
                    sel_badvaddr? badvaddr : 32'd0;

// �жϼ���߼�
// �ж����������жϹ��� && ��Ӧ�ж�ʹ�� && ȫ���ж�ʹ�� && �����쳣����
assign c0_int = |(cause_ip[7:0] & status_im[7:0]) & status_ie & !status_exl;

// �쳣/���ض����źţ������жϣ�
// ע�⣺�����쳣������syscall/break����ͨ��ex_valid_i���ݣ���������ֻ��Ҫ���ex_valid_i
assign cancel    = (ex_valid_i | eret | c0_int) && wb_over;
assign exc_valid = (ex_valid_i | eret | c0_int) && wb_valid;
assign exc_pc    = eret ? epc : `EXC_ENTER_ADDR;

endmodule
