`timescale 1ns / 1ps
//*************************************************************************
//   > �ļ���: pipeline_cpu.v
//   > ����  :�弶��ˮCPUģ�飬��ʵ��XX��ָ��
//   >        ָ��rom������ram��ʵ����xilinx IP�õ���Ϊͬ����д
//   > ����  : LOONGSON
//   > ����  : 2016-04-14
//*************************************************************************

`define IF_ID_BUS_WIDTH     64
`define ID_EXE_BUS_WIDTH    168
`define EXE_MEM_BUS_WIDTH   155
`define MEM_WB_BUS_WIDTH    156
`define JBR_BUS_WIDTH       33
`define EXC_BUS_WIDTH       33


module pipeline_cpu(
    input clk,
    input resetn,

    // display
    input  [4:0] rf_addr,
    output [31:0] rf_data,
    output [31:0] IF_pc,
    output [31:0] IF_inst,
    output [31:0] ID_pc,
    output [31:0] EXE_pc,
    output [31:0] MEM_pc,
    output [31:0] WB_pc,

    // debug
    output [31:0] cpu_5_valid,
    output [31:0] HI_data,
    output [31:0] LO_data,
    output [31:0] CP0_STATUS,
    output [31:0] CP0_CAUSE,
    output [31:0] CP0_EPC,

    //==================================================
    // AXI MASTER (INSTR)
    //==================================================
    output [31:0] M_AXI_INSTR_AWADDR,
    output [7:0]  M_AXI_INSTR_AWLEN,
    output        M_AXI_INSTR_AWVALID,
    input         M_AXI_INSTR_AWREADY,

    output [31:0] M_AXI_INSTR_WDATA,
    output        M_AXI_INSTR_WVALID,
    output        M_AXI_INSTR_WLAST,
    input         M_AXI_INSTR_WREADY,

    input  [1:0]  M_AXI_INSTR_BRESP,
    input         M_AXI_INSTR_BVALID,
    output        M_AXI_INSTR_BREADY,

    output [31:0] M_AXI_INSTR_ARADDR,
    output [7:0]  M_AXI_INSTR_ARLEN,
    output        M_AXI_INSTR_ARVALID,
    input         M_AXI_INSTR_ARREADY,

    input  [31:0] M_AXI_INSTR_RDATA,
    input         M_AXI_INSTR_RLAST,
    input         M_AXI_INSTR_RVALID,
    output        M_AXI_INSTR_RREADY,

    output [2:0]  M_AXI_INSTR_AWSIZE,
    output [2:0]  M_AXI_INSTR_ARSIZE,

    //==================================================
    // AXI MASTER (DATA)
    //==================================================
    output [31:0] M_AXI_DATA_AWADDR,
    output [7:0]  M_AXI_DATA_AWLEN,
    output        M_AXI_DATA_AWVALID,
    input         M_AXI_DATA_AWREADY,

    output [31:0] M_AXI_DATA_WDATA,
    output        M_AXI_DATA_WVALID,
    output        M_AXI_DATA_WLAST,
    input         M_AXI_DATA_WREADY,

    input  [1:0]  M_AXI_DATA_BRESP,
    input         M_AXI_DATA_BVALID,
    output        M_AXI_DATA_BREADY,

    output [31:0] M_AXI_DATA_ARADDR,
    output [7:0]  M_AXI_DATA_ARLEN,
    output        M_AXI_DATA_ARVALID,
    input         M_AXI_DATA_ARREADY,

    input  [31:0] M_AXI_DATA_RDATA,
    input         M_AXI_DATA_RLAST,
    input         M_AXI_DATA_RVALID,
    output        M_AXI_DATA_RREADY,

    output [2:0]  M_AXI_DATA_AWSIZE,
    output [2:0]  M_AXI_DATA_ARSIZE
);

// FETCH AXI user signals
wire        fetch_axi_start;
// wire [31:0] fetch_addr;
wire [31:0] fetch_axi_addr;


// MEM AXI user signals
wire        mem_axi_start;
wire        mem_axi_rw;       // 1=load, 0=store
wire [31:0] mem_axi_addr;
wire [31:0] mem_axi_wdata;
wire [7:0]  mem_axi_len;
wire        mem_axi_wvalid;
wire        mem_axi_wready;
// debug for data AXI
always @(posedge clk) begin
    if (mem_axi_start) begin
        $display("PIPE_AXI_DATA: start rw=%b addr=%h len=%0d", mem_axi_rw, mem_axi_addr, mem_axi_len);
    end
end
// --------------------------------
// AXI MASTER FOR INSTRUCTION FETCH
//-------------------------------------------------------
wire instr_user_busy;
wire instr_user_done;
wire instr_user_rvalid;
wire [31:0] instr_user_rdata;

axi_full_master #(
    .C_M_TARGET_SLAVE_BASE_ADDR(32'h00000000)
) U_AXI_INSTR (
    .M_AXI_ACLK(clk),
    .M_AXI_ARESETN(resetn),

    // AXI �������
    .M_AXI_AWID(),
    .M_AXI_AWADDR(M_AXI_INSTR_AWADDR),
    .M_AXI_AWLEN (M_AXI_INSTR_AWLEN),
    // .M_AXI_AWSIZE(),
    // .M_AXI_AWBURST(),
    .M_AXI_AWLOCK(),
    .M_AXI_AWCACHE(),
    .M_AXI_AWPROT(),
    .M_AXI_AWQOS(),
    .M_AXI_AWUSER(),
    .M_AXI_AWVALID(M_AXI_INSTR_AWVALID),
    .M_AXI_AWREADY(M_AXI_INSTR_AWREADY),

    .M_AXI_AWSIZE(M_AXI_INSTR_AWSIZE),
    .M_AXI_ARSIZE(M_AXI_INSTR_ARSIZE),

    .M_AXI_WDATA(M_AXI_INSTR_WDATA),
    .M_AXI_WSTRB(),
    .M_AXI_WLAST(M_AXI_INSTR_WLAST),
    .M_AXI_WUSER(),
    .M_AXI_WVALID(M_AXI_INSTR_WVALID),
    .M_AXI_WREADY(M_AXI_INSTR_WREADY),

    .M_AXI_BID(),
    .M_AXI_BRESP(M_AXI_INSTR_BRESP),
    .M_AXI_BUSER(),
    .M_AXI_BVALID(M_AXI_INSTR_BVALID),
    .M_AXI_BREADY(M_AXI_INSTR_BREADY),

    .M_AXI_ARID(),
    .M_AXI_ARADDR(M_AXI_INSTR_ARADDR),
    .M_AXI_ARLEN (M_AXI_INSTR_ARLEN),
    // .M_AXI_ARSIZE(),
    // .M_AXI_ARBURST(),
    .M_AXI_ARLOCK(),
    .M_AXI_ARCACHE(),
    .M_AXI_ARPROT(),
    .M_AXI_ARQOS(),
    .M_AXI_ARUSER(),
    .M_AXI_ARVALID(M_AXI_INSTR_ARVALID),
    .M_AXI_ARREADY(M_AXI_INSTR_ARREADY),

    .M_AXI_RID(),
    .M_AXI_RDATA(M_AXI_INSTR_RDATA),
    .M_AXI_RRESP(),
    .M_AXI_RLAST(M_AXI_INSTR_RLAST),
    .M_AXI_RUSER(),
    .M_AXI_RVALID(M_AXI_INSTR_RVALID),
    .M_AXI_RREADY(M_AXI_INSTR_RREADY),

    //---------------------------------------------------
    // USER ���ƽӿڣ�Fetch ʹ�ã�
    //---------------------------------------------------
    .user_start   (fetch_axi_start), 
    .user_rw      (1'b1),            // �̶�Ϊ read
    .user_addr(fetch_axi_addr),      // fetch.v �е� PC
    .user_len     (8'd1),            // ÿ�ζ�1��ָ��

    .user_wdata   (32'd0),           // �����õ�
    .user_wvalid  (1'b0),
    .user_wready  (),

    .user_rdata   (instr_user_rdata),
    .user_rvalid  (instr_user_rvalid),
    .user_rready  (1'b1),

    .user_busy    (instr_user_busy),
    .user_done    (instr_user_done),
    .user_error   ()
);

//-------------------------------------------------------
// AXI MASTER FOR DATA LOAD/STORE
//-------------------------------------------------------
wire data_user_busy;
wire data_user_done;
wire [31:0] data_user_rdata;
wire data_user_rvalid;

axi_full_master #(
    .C_M_TARGET_SLAVE_BASE_ADDR(32'h00000000)
) U_AXI_DATA (
    .M_AXI_ACLK(clk),
    .M_AXI_ARESETN(resetn),

    // AXI �������
    .M_AXI_AWID(),
    .M_AXI_AWADDR(M_AXI_DATA_AWADDR),
    .M_AXI_AWLEN (M_AXI_DATA_AWLEN),
    // .M_AXI_AWSIZE(),
    // .M_AXI_AWBURST(),
    .M_AXI_AWLOCK(),
    .M_AXI_AWCACHE(),
    .M_AXI_AWPROT(),
    .M_AXI_AWQOS(),
    .M_AXI_AWUSER(),
    .M_AXI_AWVALID(M_AXI_DATA_AWVALID),
    .M_AXI_AWREADY(M_AXI_DATA_AWREADY),

    .M_AXI_AWSIZE(M_AXI_DATA_AWSIZE),
    .M_AXI_ARSIZE(M_AXI_DATA_ARSIZE),

    .M_AXI_WDATA(M_AXI_DATA_WDATA),
    .M_AXI_WSTRB(),
    .M_AXI_WLAST(M_AXI_DATA_WLAST),
    .M_AXI_WUSER(),
    .M_AXI_WVALID(M_AXI_DATA_WVALID),
    .M_AXI_WREADY(M_AXI_DATA_WREADY),

    .M_AXI_BID(),
    .M_AXI_BRESP(M_AXI_DATA_BRESP),
    .M_AXI_BUSER(),
    .M_AXI_BVALID(M_AXI_DATA_BVALID),
    .M_AXI_BREADY(M_AXI_DATA_BREADY),

    .M_AXI_ARID(),
    .M_AXI_ARADDR(M_AXI_DATA_ARADDR),
    .M_AXI_ARLEN (M_AXI_DATA_ARLEN),
    // .M_AXI_ARSIZE(),
    // .M_AXI_ARBURST(),
    .M_AXI_ARLOCK(),
    .M_AXI_ARCACHE(),
    .M_AXI_ARPROT(),
    .M_AXI_ARQOS(),
    .M_AXI_ARUSER(),
    .M_AXI_ARVALID(M_AXI_DATA_ARVALID),
    .M_AXI_ARREADY(M_AXI_DATA_ARREADY),

    .M_AXI_RID(),
    .M_AXI_RDATA(M_AXI_DATA_RDATA),
    .M_AXI_RRESP(),
    .M_AXI_RLAST(M_AXI_DATA_RLAST),
    .M_AXI_RUSER(),
    .M_AXI_RVALID(M_AXI_DATA_RVALID),
    .M_AXI_RREADY(M_AXI_DATA_RREADY),

    //---------------------------------------------------
    // USER �ӿ� (mem ʹ��)
    //---------------------------------------------------
    .user_start   (mem_axi_start),
    .user_rw      (mem_axi_rw),        // 0 = store, 1 = load
    .user_addr    (mem_axi_addr),
    .user_len     (mem_axi_len),

    .user_wdata   (mem_axi_wdata),
    .user_wvalid  (mem_axi_wvalid),
    .user_wready  (mem_axi_wready),

    .user_rdata   (data_user_rdata),
    .user_rvalid  (data_user_rvalid),
    .user_rready  (1'b1),

    .user_busy    (data_user_busy),
    .user_done    (data_user_done),
    .user_error   ()
);



//------------------------{5����ˮ�����ź�}begin-------------------------//
    //5ģ���valid�ź�
    reg IF_valid;
    reg ID_valid;
    reg EXE_valid;
    reg MEM_valid;
    reg WB_valid;
    //5ģ��ִ������ź�,���Ը�ģ������
    wire IF_over;
    wire ID_over;
    wire EXE_over;
    wire MEM_over;
    wire WB_over;
    //5ģ��������һ��ָ�����
    wire IF_allow_in;
    wire ID_allow_in;
    wire EXE_allow_in;
    wire MEM_allow_in;
    wire WB_allow_in;
    
    // syscall��eret����д�ؼ�ʱ�ᷢ��cancel�źţ�
    wire cancel;    // ȡ���Ѿ�ȡ��������������ˮ��ִ�е�ָ��
    
    //������������ź�:������Ч���򱾼�ִ��������¼��������
    assign IF_allow_in  = (IF_over & ID_allow_in) | cancel;
    assign ID_allow_in  = ~ID_valid  | (ID_over  & EXE_allow_in);
    assign EXE_allow_in = ~EXE_valid | (EXE_over & MEM_allow_in);
    assign MEM_allow_in = ~MEM_valid | (MEM_over & WB_allow_in );
    assign WB_allow_in  = ~WB_valid  | WB_over;
   
    //IF_valid���ڸ�λ��һֱ��Ч
   always @(posedge clk)
    begin
        if (!resetn)
        begin
            IF_valid <= 1'b0;
        end
        else
        begin
            IF_valid <= 1'b1;
        end
    end
    
    //ID_valid
    always @(posedge clk)
    begin
        if (!resetn || cancel)
        begin
            ID_valid <= 1'b0;
        end
        else if (ID_allow_in)
        begin
            ID_valid <= IF_over;
        end
    end
    
    //EXE_valid
    always @(posedge clk)
    begin
        if (!resetn || cancel)
        begin
            EXE_valid <= 1'b0;
        end
        else if (EXE_allow_in)
        begin
            EXE_valid <= ID_over;
        end
    end
    
    //MEM_valid
    always @(posedge clk)
    begin
        if (!resetn || cancel)
        begin
            MEM_valid <= 1'b0;
        end
        else if (MEM_allow_in)
        begin
            MEM_valid <= EXE_over;
        end
    end
    
    //WB_valid
    always @(posedge clk)
    begin
        if (!resetn || cancel)
        begin
            WB_valid <= 1'b0;
        end
        else if (WB_allow_in)
        begin
            WB_valid <= MEM_over;
        end
    end
    
    //չʾ5����valid�ź�
    assign cpu_5_valid = {12'd0         ,{4{IF_valid }},{4{ID_valid}},
                          {4{EXE_valid}},{4{MEM_valid}},{4{WB_valid}}};
//-------------------------{5����ˮ�����ź�}end--------------------------//

//--------------------------{5���������}begin---------------------------//
    wire [ 63:0] IF_ID_bus;   // IF->ID������
    wire [167:0] ID_EXE_bus;  // ID->EXE������
    wire [154:0] EXE_MEM_bus; // EXE->MEM������
    wire [155:0] MEM_WB_bus;  // MEM->WB������
    
    //�������������ź�
    reg [ 63:0] IF_ID_bus_r;
    reg [167:0] ID_EXE_bus_r;
    reg [154:0] EXE_MEM_bus_r;
    reg [155:0] MEM_WB_bus_r;
    
    //IF��ID�������ź�
    always @(posedge clk)
    begin
        if(IF_over && ID_allow_in)
        begin
            IF_ID_bus_r <= IF_ID_bus;
        end
    end
    //ID��EXE�������ź�
    always @(posedge clk)
    begin
        if(ID_over && EXE_allow_in)
        begin
            ID_EXE_bus_r <= ID_EXE_bus;
        end
    end
    //EXE��MEM�������ź�
    always @(posedge clk)
    begin
        if(EXE_over && MEM_allow_in)
        begin
            EXE_MEM_bus_r <= EXE_MEM_bus;
        end
    end    
    //MEM��WB�������ź�
    always @(posedge clk)
    begin
        if(MEM_over && WB_allow_in)
        begin
            MEM_WB_bus_r <= MEM_WB_bus;
        end
    end
//---------------------------{5���������}end----------------------------//

//------------------------{��·����ź�}begin---------------------------//

    // ��·�����ź�
    wire [31:0] EXE_result;    // EXE�����
    wire [31:0] MEM_result;    // MEM�����  
    wire [31:0] WB_result;     // WB�����
    
    // ��·�����ź�
    wire [4:0] EXE_wdest;      // EXE��д��Ŀ��Ĵ���
    wire [4:0] MEM_wdest;      // MEM��д��Ŀ��Ĵ���
    wire [4:0] WB_wdest;       // WB��д��Ŀ��Ĵ���
    
    // EXE��ָ��������Ϣ
    wire EXE_inst_load;        // EXE��Loadָ��
    wire EXE_inst_mult;        // EXE���˷�ָ��
    
//------------------------{��·����ź�}end----------------------------//

//--------------------------{���������ź�}begin--------------------------//
    //��ת����
    wire [ 32:0] jbr_bus;    

    //IF��inst_rom����
    // wire [31:0] inst_addr;
    // wire [31:0] inst;

    //ID��EXE��MEM��WB����
    wire [ 4:0] EXE_wdest;
    wire [ 4:0] MEM_wdest;
    wire [ 4:0] WB_wdest;
    
    //MEM��data_ram����    
    // wire [ 3:0] dm_wen;
    // wire [31:0] dm_addr;
    // wire [31:0] dm_wdata;
    // wire [31:0] dm_rdata;

    //ID��regfile����
    wire [ 4:0] rs;
    wire [ 4:0] rt;   
    wire [31:0] rs_value;
    wire [31:0] rt_value;
    
    //WB��regfile����
    wire        rf_wen;
    wire [ 4:0] rf_wdest;
    wire [31:0] rf_wdata;    
    
    //WB��IF��Ľ����ź�
    wire [ 32:0] exc_bus;
//---------------------------{���������ź�}end---------------------------//

//-------------------------{��ģ��ʵ����}begin---------------------------//
    wire next_fetch; //��������ȡָģ�飬��Ҫ������PCֵ
    //IF�������ʱ��������PCֵ��ȡ��һ��ָ��
    assign next_fetch = IF_allow_in;
    fetch IF_module(             // ȡָ��
        .clk       (clk       ),  // I, 1
        .resetn    (resetn    ),  // I, 1
        .IF_valid  (IF_valid  ),  // I, 1
        .next_fetch(next_fetch),  // I, 1
        // .inst      (inst      ),  // I, 32
        .jbr_bus   (jbr_bus   ),  // I, 33
        // .inst_addr (inst_addr ),  // O, 32
        .IF_over   (IF_over   ),  // O, 1
        .IF_ID_bus (IF_ID_bus ),  // O, 64

        .axi_start   (fetch_axi_start),
        .axi_done    (instr_user_done),
        .axi_rdata   (instr_user_rdata),
        .axi_busy    (instr_user_busy),
        .axi_addr(fetch_axi_addr),
        
        //5����ˮ�����ӿ�
        .exc_bus   (exc_bus   ),  // I, 32
        
        //չʾPC��ȡ����ָ��
        .IF_pc     (IF_pc     ),  // O, 32
        .IF_inst   (IF_inst   )   // O, 32
    );

    // inst = axi_rdata;
    // IF_over = axi_done;

    decode ID_module(               // ���뼶
        .clk        (clk        ),  // I, 1
        .ID_valid   (ID_valid   ),  // I, 1
        .IF_ID_bus_r(IF_ID_bus_r),  // I, 64
        .rs_value   (rs_value   ),  // I, 32
        .rt_value   (rt_value   ),  // I, 32
        .rs         (rs         ),  // O, 5
        .rt         (rt         ),  // O, 5
        .jbr_bus    (jbr_bus    ),  // O, 33
//        .inst_jbr   (inst_jbr   ),  // O, 1
        .ID_over    (ID_over    ),  // O, 1
        .ID_EXE_bus (ID_EXE_bus ),  // O, 167
        
        //5����ˮ����
        .IF_over     (IF_over     ),// I, 1
        .EXE_wdest   (EXE_wdest   ),// I, 5
        .MEM_wdest   (MEM_wdest   ),// I, 5
        .WB_wdest    (WB_wdest    ),// I, 5

        // ��·��
        .EXE_result(EXE_result),  // I, 32
        .MEM_result(MEM_result),  // I, 32
        .WB_result(WB_result),    // I, 32

        .EXE_valid(EXE_valid),    // I, 1
        .MEM_valid(MEM_valid),    // I, 1
        .WB_valid(WB_valid),      // I, 1
        
        // EXE��ָ��������Ϣ
        .EXE_inst_load(EXE_inst_load),  // I, 1
        .EXE_inst_mult(EXE_inst_mult),  // I, 1
        
        //չʾPC
        .ID_pc       (ID_pc       ) // O, 32
    ); 

    exe EXE_module(                   // ִ�м�
        .EXE_valid   (EXE_valid   ),  // I, 1
        .ID_EXE_bus_r(ID_EXE_bus_r),  // I, 167
        .EXE_over    (EXE_over    ),  // O, 1 
        .EXE_MEM_bus (EXE_MEM_bus ),  // O, 154
        
        //5����ˮ����
        .clk         (clk         ),  // I, 1
        .EXE_wdest   (EXE_wdest   ),  // O, 5

        // ��·��������
        .EXE_result(EXE_result),  // O, 32
        
        // EXE��ָ��������Ϣ���
        .EXE_inst_load(EXE_inst_load),  // O, 1
        .EXE_inst_mult(EXE_inst_mult),  // O, 1
        
        //չʾPC
        .EXE_pc      (EXE_pc      )   // O, 32
    );

    mem MEM_module(                     // �ô漶
        .clk          (clk          ),  // I, 1 
        .MEM_valid    (MEM_valid    ),  // I, 1
        .EXE_MEM_bus_r(EXE_MEM_bus_r),  // I, 155
        // .dm_rdata     (dm_rdata     ),  // I, 32
        // .dm_addr      (dm_addr      ),  // O, 32
        // .dm_wen       (dm_wen       ),  // O, 4 
        // .dm_wdata     (dm_wdata     ),  // O, 32
        .MEM_over     (MEM_over     ),  // O, 1
        .MEM_WB_bus   (MEM_WB_bus   ),  // O, 156
        
        //5����ˮ�����ӿ�
        .MEM_allow_in (MEM_allow_in ),  // I, 1
        .MEM_wdest    (MEM_wdest    ),  // O, 5

        // ������·�������
        .MEM_result(MEM_result),  // O, 32
        
        .axi_start   (mem_axi_start),
        .axi_rw      (mem_axi_rw),
        .axi_addr    (mem_axi_addr),
        .axi_len     (mem_axi_len),
        .axi_wdata   (mem_axi_wdata),

        .axi_rdata   (data_user_rdata),
        .axi_rvalid  (data_user_rvalid),
        .axi_done    (data_user_done),
        .axi_busy    (data_user_busy),
        .axi_wvalid  (mem_axi_wvalid),
        .axi_wready  (mem_axi_wready),

        //չʾPC
        .MEM_pc       (MEM_pc       )   // O, 32
    );          
 
    wb WB_module(                     // д�ؼ�
        .WB_valid    (WB_valid    ),  // I, 1
        .MEM_WB_bus_r(MEM_WB_bus_r),  // I, 156
        .rf_wen      (rf_wen      ),  // O, 1
        .rf_wdest    (rf_wdest    ),  // O, 5
        .rf_wdata    (rf_wdata    ),  // O, 32
          .WB_over     (WB_over     ),  // O, 1
        
        //5����ˮ�����ӿ�
        .clk         (clk         ),  // I, 1
      .resetn      (resetn      ),  // I, 1
        .exc_bus     (exc_bus     ),  // O, 32
        .WB_wdest    (WB_wdest    ),  // O, 5
        .cancel      (cancel      ),  // O, 1
        
        // ������·�������
        .WB_result(WB_result),  // O, 32
        
        //չʾPC��HI/LOֵ
        .WB_pc       (WB_pc       ),  // O, 32
        .HI_data     (HI_data     ),  // O, 32
        .LO_data     (LO_data     ),  // O, 32
        // ����CP0�Ĵ���
        .cp0_status  (CP0_STATUS  ),  // O, 32
        .cp0_cause   (CP0_CAUSE   ),  // O, 32
        .cp0_epc     (CP0_EPC     )   // O, 32
    );

    // inst_rom inst_rom_module(         // ָ��洢��
    //     .clka       (clk           ),  // I, 1 ,ʱ��
    //     .addra      (inst_addr[9:2]),  // I, 8 ,ָ���ַ
    //     .douta      (inst          )   // O, 32,ָ��
    // );

    regfile rf_module(        // �Ĵ�����ģ��
        .clk    (clk      ),  // I, 1
        .wen    (rf_wen   ),  // I, 1
        .raddr1 (rs       ),  // I, 5
        .raddr2 (rt       ),  // I, 5
        .waddr  (rf_wdest ),  // I, 5
        .wdata  (rf_wdata ),  // I, 32
        .rdata1 (rs_value ),  // O, 32
        .rdata2 (rt_value ),  // O, 32

        //display rf
        .test_addr(rf_addr),  // I, 5
        .test_data(rf_data)   // O, 32
    );
    
    // data_ram data_ram_module(   // ���ݴ洢ģ��
    //     .clka   (clk         ),  // I, 1,  ʱ��
    //     .wea    (dm_wen      ),  // I, 1,  дʹ��
    //     .addra  (dm_addr[9:2]),  // I, 8,  ����ַ
    //     .dina   (dm_wdata    ),  // I, 32, д����
    //     .douta  (dm_rdata    ),  // O, 32, ������

    //     //display mem
    //     .clkb   (clk          ),  // I, 1,  ʱ��
    //     .web    (4'd0         ),  // ��ʹ�ö˿�2��д����
    //     .addrb  (mem_addr[9:2]),  // I, 8,  ����ַ
    //     .doutb  (mem_data     ),  // I, 32, д����
    //     .dinb   (32'd0        )   // ��ʹ�ö˿�2��д����
    // );
//--------------------------{��ģ��ʵ����}end----------------------------//
endmodule
