`timescale 1ns / 1ps
`define STARTADDR 32'H00000000

module fetch(
    input             clk,
    input             resetn,
    input             IF_valid,
    input             next_fetch,      // pipeline �������
    input      [32:0] jbr_bus,        // ��ת����

    // ===== AXI USER INTERFACE =====
    output reg        axi_start,      // ���� 1 ���ڿ�ʼ AXI read
    output reg [31:0] axi_addr,       // AXI ����ַ (PC)
    input             axi_done,       // AXI ������� = inst ��Ч
    input      [31:0] axi_rdata,      // AXI ������ָ��
    input             axi_busy,       // AXI ����ִ��

    //===============================
    // pipeline ���
    //===============================
    output reg        IF_over,        // ���
    output     [63:0] IF_ID_bus,      // {PC , INST}

    // �쳣
    input      [32:0] exc_bus,

    // debug
    output     [31:0] IF_pc,
    output     [31:0] IF_inst
);

    //===================== PC �߼� =======================
    reg  [31:0] pc;
    reg  [31:0] inst_reg;   // ��ָ���һ�ı��棬���� AXI ���߿���ʱ�� 0

    wire [31:0] next_pc;
    wire [31:0] seq_pc;

    // ��ת
    wire        jbr_taken;
    wire [31:0] jbr_target;
    assign {jbr_taken, jbr_target} = jbr_bus;

    // �쳣
    wire        exc_valid;
    wire [31:0] exc_pc;
    assign {exc_valid, exc_pc} = exc_bus;

    // PC + 4
    assign seq_pc = pc + 32'd4;

    // PC ѡ��
    assign next_pc = exc_valid ? exc_pc :
                     jbr_taken ? jbr_target :
                     seq_pc;

    // **ע�⣺ֻ�е�ǰָ������"ȡ�ز��ұ���ˮ����"ʱ�Ÿ��� PC**
    always @(posedge clk) begin
        if (!resetn)
            pc <= `STARTADDR;
        // ֻ�С���һ��ָ����ȡ��(=IF_over)������ˮ���������(next_fetch)
        // ʱ�Ÿ��� PC������ axi_done ������ next_fetch ��λ���� PC ��ס
        else if (next_fetch && IF_over)
            pc <= next_pc;
    end

    // ָ���һ�ı��棨AXI ���߿���ʱ IF_inst ����������
    always @(posedge clk) begin
        if (!resetn)
            inst_reg <= 32'h0;
        else if (axi_done)
            inst_reg <= axi_rdata;
    end

    //===================== AXI �����񴥷� ======================
    // ʹ�ô�ͳparameter����״̬��
    parameter [1:0] IDLE = 2'b00,
                  REQUEST = 2'b01,
                  PENDING = 2'b10,
                  DONE = 2'b11;

    reg [1:0] current_state, next_state;

    always @(posedge clk) begin
        if (!resetn)
            current_state <= IDLE;
        else
            current_state <= next_state;
    end

    always @(*) begin
        case(current_state)
            IDLE: begin
                if (IF_valid && !axi_busy)
                    next_state = REQUEST;
                else
                    next_state = IDLE;
            end
            REQUEST: begin
                next_state = PENDING;  // �����������������PENDING״̬
            end
            PENDING: begin
                if (axi_done)
                    next_state = DONE;
                else
                    next_state = PENDING;
            end
            DONE: begin
                if (next_fetch)
                    next_state = IDLE;
                else
                    next_state = DONE;
            end
            default: next_state = IDLE;
        endcase
    end

    // AXI �����ź�
    always @(posedge clk) begin
        if (!resetn) begin
            axi_start <= 1'b0;
            axi_addr  <= `STARTADDR;
        end
        else begin
            // �� REQUEST ״̬���� 1 �����壬�����浱ǰ PC Ϊ AXI ��ַ
            axi_start <= (current_state == REQUEST);
            if (current_state == REQUEST) begin
                axi_addr <= pc;
                $display("Time=%0t FETCH: Requesting PC=%h", $time, pc);
            end
        end
    end

    //===================== IF_over ���� ======================
    // IF_over ��Ϊ���ֻ��ƣ�axi_done ��λ��next_fetch ���ͱ�ʾ�¼��ѽ���
    always @(posedge clk) begin
        if (!resetn)
            IF_over <= 1'b0;
        else if (axi_done)
            IF_over <= 1'b1;          // ָ����ȡ��
        else if (next_fetch)
            IF_over <= 1'b0;          // �¼��ѽ��գ�׼����һ��
    end

    //===================== ��� ======================
    assign IF_ID_bus = { pc, inst_reg };
    assign IF_pc     = pc;
    assign IF_inst   = inst_reg;   // �ô��ĺ�� inst_reg�����β������Ǳ� 0

endmodule