`timescale 1ns / 1ps
`define STARTADDR 32'H00000034

module fetch(
    input             clk,
    input             resetn,
    input             IF_valid,
    input             next_fetch,      // pipeline �������
    input      [32:0] jbr_bus,        // ��ת����

    // ===== AXI USER INTERFACE =====
    output reg        axi_start,      // ���� 1 ���ڿ�ʼ AXI read
    output reg [31:0] axi_addr,       // AXI ����ַ (PC)
    input             axi_done,       // AXI ������� = inst ��Ч
    input      [31:0] axi_rdata,      // AXI ������ָ��
    input             axi_busy,       // AXI ����ִ��

    //===============================
    // pipeline ���
    //===============================
    output reg        IF_over,        // ���
    output     [63:0] IF_ID_bus,      // {PC , INST}

    // �쳣
    input      [32:0] exc_bus,

    // debug
    output     [31:0] IF_pc,
    output     [31:0] IF_inst
);

    //===================== PC �߼� =======================
    reg  [31:0] pc;
    reg  [31:0] inst_reg;   // ��ָ���һ�ı��棬���� AXI ���߿���ʱ�� 0

    wire [31:0] next_pc;
    wire [31:0] seq_pc;

    // ��ת
    wire        jbr_taken;
    wire [31:0] jbr_target;
    assign {jbr_taken, jbr_target} = jbr_bus;

    // �쳣
    wire        exc_valid;
    wire [31:0] exc_pc;
    assign {exc_valid, exc_pc} = exc_bus;

    // PC + 4
    assign seq_pc = { pc[31:2] + 1'b1, pc[1:0] };

    // PC ѡ��
    assign next_pc = exc_valid ? exc_pc :
                     jbr_taken ? jbr_target :
                     seq_pc;

    // **ע�⣺ֻ�е�ǰָ��������ȡ�ز��ұ���ˮ���ܡ�ʱ�Ÿ��� PC**
    always @(posedge clk) begin
        if (!resetn)
            pc <= `STARTADDR;
        else if (next_fetch && axi_done)
            pc <= next_pc;
    end

    // ָ���һ�ı��棨AXI ���߿���ʱ IF_inst ����������
    always @(posedge clk) begin
        if (!resetn)
            inst_reg <= 32'h0;
        else if (axi_done)
            inst_reg <= axi_rdata;
    end

    //===================== AXI �����񴥷� ======================
    // �ǳ��򵥵�״̬������֤����ʱ�����ֻ���� 1 ��������
    reg started;        // �Ƿ��Ѿ�������һ�ζ�
    reg outstanding;    // �Ƿ��ж��������ڽ�����

    always @(posedge clk) begin
        if (!resetn) begin
            axi_start   <= 1'b0;
            axi_addr    <= `STARTADDR;
            started     <= 1'b0;
            outstanding <= 1'b0;
        end
        else begin
            axi_start <= 1'b0;   // Ĭ������

            // ��ǰָ�������
            if (axi_done)
                outstanding <= 1'b0;

            // ��λ���һ�Σ�ֱ�Ӱ���ǰ pc ȡһ��ָ��
            if (!started && !outstanding && !axi_busy) begin
                axi_start   <= 1'b1;
                axi_addr    <= pc;         // ������ STARTADDR
                started     <= 1'b1;
                outstanding <= 1'b1;
            end
            // ��������ǰû�й�������ʱ����ȡ��һ��ָ��
            else if (started && !outstanding && !axi_busy && IF_valid) begin
                axi_start   <= 1'b1;
                axi_addr    <= pc;         // ע�⣺pc �Ѿ�����һ�� axi_done ʱ����Ϊ��һ��
                outstanding <= 1'b1;
            end
        end
    end

    //===================== IF_over ���� ======================
    // AXI ����� -> IF �����
    always @(posedge clk) begin
        if (!resetn)
            IF_over <= 1'b0;
        else
            IF_over <= axi_done;
    end

    //===================== ��� ======================
    assign IF_ID_bus = { pc, inst_reg };
    assign IF_pc     = pc;
    assign IF_inst   = inst_reg;   // �ô��ĺ�� inst_reg�����β������Ǳ� 0

endmodule
